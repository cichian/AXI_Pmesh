module test(

);

`ifdef TEST
    $display ("test");
`else 
    $display ("no test");
`endif





endmodule